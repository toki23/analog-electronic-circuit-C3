* Rc直列回路
V 1 0 sin(0V 1V 50Hz)
R 2 0 1k
C 1 2 1u 
.tran 0.1ms 40ms 20ms
.control
    run
    plot v(1),v(2)
.endc
.end